module contagemRegressiva(
    input umSegundo,
    input aspersao,
    input gotejamento,
    input casoEspecifico,
    input [2:0] nivelDagua,
    input button,
    output [3:0] Us, Ds, Um, Dm
);

endmodule
